`define A 1
